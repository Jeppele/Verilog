module counter #(
    parameter N = 10
) (
    port_list
);
    
endmodule